   
    parameter PROC_NUM = 11;
    parameter ST_IDLE = 3'b000;
    parameter ST_FILTER_FAKE = 3'b001;
    parameter ST_DL_DETECTED = 3'b010;
    parameter ST_DL_REPORT = 3'b100;
   

    reg [2:0] CS_fsm;
    reg [2:0] NS_fsm;
    reg [PROC_NUM - 1:0] dl_detect_reg;
    reg [PROC_NUM - 1:0] dl_done_reg;
    reg [PROC_NUM - 1:0] origin_reg;
    reg [PROC_NUM - 1:0] dl_in_vec_reg;
    reg [31:0] dl_keep_cnt;
    reg stop_report_path;
    reg [PROC_NUM - 1:0] reported_proc;
    integer i;
    integer fp;

    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            reported_proc <= 'b0;
        end
        else if (CS_fsm == ST_DL_REPORT) begin
            reported_proc <= reported_proc | dl_in_vec;
        end
        else if (CS_fsm == ST_DL_DETECTED) begin
            reported_proc <= 'b0;
        end
    end

    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            stop_report_path <= 1'b0;
        end
        else if (CS_fsm == ST_DL_REPORT && (|(dl_in_vec & reported_proc))) begin
            stop_report_path <= 1'b1;
        end
        else if (CS_fsm == ST_IDLE) begin
            stop_report_path <= 1'b0;
        end
    end

    // FSM State machine
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            CS_fsm <= ST_IDLE;
        end
        else begin
            CS_fsm <= NS_fsm;
        end
    end

    always @ (CS_fsm or dl_in_vec or dl_detect_reg or dl_done_reg or dl_in_vec or origin_reg or dl_keep_cnt) begin
        case (CS_fsm)
            ST_IDLE : begin
                if (|dl_in_vec) begin
                    NS_fsm = ST_FILTER_FAKE;
                end
                else begin
                    NS_fsm = ST_IDLE;
                end
            end
            ST_FILTER_FAKE: begin
                if (dl_keep_cnt >= 32'd1000) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else if (dl_detect_reg != (dl_detect_reg & dl_in_vec)) begin
                    NS_fsm = ST_IDLE;
                end
                else begin
                    NS_fsm = ST_FILTER_FAKE;
                end
            end
            ST_DL_DETECTED: begin
                // has unreported deadlock cycle
                if ((dl_detect_reg != dl_done_reg) && stop_report_path == 1'b0) begin
                    NS_fsm = ST_DL_REPORT;
                end
                else begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
            ST_DL_REPORT: begin
                if (|(dl_in_vec & origin_reg)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                // avoid report deadlock ring.
                else if (|(dl_in_vec & reported_proc)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else begin
                    NS_fsm = ST_DL_REPORT;
                end
            end
            default: NS_fsm = ST_IDLE;
        endcase
    end

    // dl_detect_reg record the procs that first detect deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_detect_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_IDLE) begin
                dl_detect_reg <= dl_in_vec;
            end
        end
    end

    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_keep_cnt <= 32'h0;
        end
        else begin
            if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg == (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= dl_keep_cnt + 32'h1;
            end
            else if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg != (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= 32'h0;
            end
        end
    end

    // dl_detect_out keeps in high after deadlock detected
    assign dl_detect_out = (|dl_detect_reg) && (CS_fsm == ST_DL_DETECTED || CS_fsm == ST_DL_REPORT);

    // dl_done_reg record the cycles has been reported
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_done_reg <= 'b0;
        end
        else begin
            if ((CS_fsm == ST_DL_REPORT) && (|(dl_in_vec & dl_detect_reg) == 'b1)) begin
                dl_done_reg <= dl_done_reg | dl_in_vec;
            end
        end
    end

    // clear token once a cycle is done
    assign token_clear = (CS_fsm == ST_DL_REPORT) ? ((|(dl_in_vec & origin_reg)) ? 'b1 : 'b0) : 'b0;

    // origin_reg record the current cycle start id
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            origin_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                origin_reg <= origin;
            end
        end
    end
   
    // origin will be valid for only one cycle
    wire [PROC_NUM*PROC_NUM - 1:0] origin_tmp;
    assign origin_tmp[PROC_NUM - 1:0] = (dl_detect_reg[0] & ~dl_done_reg[0]) ? 'b1 : 'b0;
    genvar j;
    generate
    for(j = 1;j < PROC_NUM;j = j + 1) begin: F1
        assign origin_tmp[j*PROC_NUM +: PROC_NUM] = (dl_detect_reg[j] & ~dl_done_reg[j]) ? ('b1 << j) : origin_tmp[(j - 1)*PROC_NUM +: PROC_NUM];
    end
    endgenerate
    always @ (CS_fsm or origin_tmp) begin
        if (CS_fsm == ST_DL_DETECTED) begin
            origin = origin_tmp[(PROC_NUM - 1)*PROC_NUM +: PROC_NUM];
        end
        else begin
            origin = 'b0;
        end
    end

    
    // dl_in_vec_reg record the current cycle dl_in_vec
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_in_vec_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                dl_in_vec_reg <= origin;
            end
            else if (CS_fsm == ST_DL_REPORT) begin
                dl_in_vec_reg <= dl_in_vec;
            end
        end
    end
    
    // find_df_deadlock to report the deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            find_df_deadlock <= 1'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED && ((dl_detect_reg == dl_done_reg) || (stop_report_path == 1'b1))) begin
                find_df_deadlock <= 1'b1;
            end
            else if (CS_fsm == ST_IDLE) begin
                find_df_deadlock <= 1'b0;
            end
        end
    end
    
    // get the first valid proc index in dl vector
    function integer proc_index(input [PROC_NUM - 1:0] dl_vec);
        begin
            proc_index = 0;
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_vec[i]) begin
                    proc_index = i;
                end
            end
        end
    endfunction

    // get the proc path based on dl vector
    function [920:0] proc_path(input [PROC_NUM - 1:0] dl_vec);
        integer index;
        begin
            index = proc_index(dl_vec);
            case (index)
                0 : begin
                    proc_path = "GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0";
                end
                1 : begin
                    proc_path = "GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0";
                end
                2 : begin
                    proc_path = "GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0";
                end
                3 : begin
                    proc_path = "GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0";
                end
                4 : begin
                    proc_path = "GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0";
                end
                5 : begin
                    proc_path = "GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0";
                end
                6 : begin
                    proc_path = "GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0";
                end
                7 : begin
                    proc_path = "GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0";
                end
                8 : begin
                    proc_path = "GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ToField_U0";
                end
                9 : begin
                    proc_path = "GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.chal2_U0";
                end
                10 : begin
                    proc_path = "GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.aggregate_coef_U0";
                end
                default : begin
                    proc_path = "unknown";
                end
            endcase
        end
    endfunction

    // print the headlines of deadlock detection
    task print_dl_head;
        begin
            $display("\n//////////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", $time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            fp = $fopen("deadlock_db.dat", "w");
        end
    endtask

    // print the start of a cycle
    task print_cycle_start(input reg [920:0] proc_path, input integer cycle_id);
        begin
            $display("/////////////////////////");
            $display("// Dependence cycle %0d:", cycle_id);
            $display("// (1): Process: %0s", proc_path);
            $fdisplay(fp, "Dependence_Cycle_ID %0d", cycle_id);
            $fdisplay(fp, "Dependence_Process_ID 1");
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print the end of deadlock detection
    task print_dl_end(input integer num, input integer record_time);
        begin
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// Totally %0d cycles detected!", num);
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", record_time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            $fdisplay(fp, "Dependence_Cycle_Number %0d", num);
            $fclose(fp);
        end
    endtask

    // print one proc component in the cycle
    task print_cycle_proc_comp(input reg [920:0] proc_path, input integer cycle_comp_id);
        begin
            $display("// (%0d): Process: %0s", cycle_comp_id, proc_path);
            $fdisplay(fp, "Dependence_Process_ID %0d", cycle_comp_id);
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print one channel component in the cycle
    task print_cycle_chan_comp(input [PROC_NUM - 1:0] dl_vec1, input [PROC_NUM - 1:0] dl_vec2);
        reg [984:0] chan_path;
        integer index1;
        integer index2;
        begin
            index1 = proc_index(dl_vec1);
            index2 = proc_index(dl_vec2);
            case (index1)
                0 : begin // for proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0'
                    case(index2)
                    2: begin //  for dep proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.k_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0.k_strm_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0.k_strm_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.k_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.k_strm_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.k_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.k_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.k_strm_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.k_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_key_to_mem_U0_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_key_to_mem_U0_U.if_full_n & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0.ap_start & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_key_to_mem_U0_U.if_read} start_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_key_to_mem_U0_U.if_full_n & grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0.ap_start & ~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_key_to_mem_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_key_to_mem_U0_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0',");
                        end
                    end
                    1: begin //  for dep proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.leaf_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0.leaf_strm_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0.leaf_strm_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.leaf_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.leaf_strm_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.leaf_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.leaf_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.leaf_strm_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.leaf_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_seed_gen_U0_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_seed_gen_U0_U.if_full_n & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0.ap_start & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_seed_gen_U0_U.if_read} start_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_seed_gen_U0_U.if_full_n & grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0.ap_start & ~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_seed_gen_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_seed_gen_U0_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0',");
                        end
                    end
                    endcase
                end
                1 : begin // for proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0'
                    case(index2)
                    0: begin //  for dep proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.leaf_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.leaf_strm_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.leaf_strm_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.leaf_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.leaf_strm_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.leaf_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.leaf_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.leaf_strm_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.leaf_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_seed_gen_U0_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_seed_gen_U0_U.if_empty_n & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.ap_idle & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_seed_gen_U0_U.if_write} start_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_seed_gen_U0_U.if_empty_n & grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.ap_idle & ~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_seed_gen_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_seed_gen_U0_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0',");
                        end
                    end
                    3: begin //  for dep proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_strm_cp_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.com_strm_cp_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.com_strm_cp_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_strm_cp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_strm_cp_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_strm_cp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_strm_cp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_strm_cp_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_strm_cp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel '' info is :
// blk sig is {{ap_done_reg_1 & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.ap_done & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0.ap_done} output_sync}
                        if ((ap_done_reg_1 & grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.ap_done & ~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0.ap_done)) begin
                            $display("//      Blocked by output sync logic with process : 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0'");
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_com_to_mem_U0_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_com_to_mem_U0_U.if_full_n & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.ap_start & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.real_start & (trans_in_cnt_1 == trans_out_cnt_1) & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_com_to_mem_U0_U.if_read} start_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_com_to_mem_U0_U.if_full_n & grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.ap_start & ~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.real_start & (trans_in_cnt_1 == trans_out_cnt_1) & ~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_com_to_mem_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_com_to_mem_U0_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0',");
                        end
                    end
                    2: begin //  for dep proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0'
// for dep channel '' info is :
// blk sig is {{ap_done_reg_1 & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.ap_done & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0.ap_done} output_sync}
                        if ((ap_done_reg_1 & grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.ap_done & ~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0.ap_done)) begin
                            $display("//      Blocked by output sync logic with process : 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0'");
                        end
                    end
                    endcase
                end
                2 : begin // for proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0'
                    case(index2)
                    0: begin //  for dep proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.k_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0.k_strm_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0.k_strm_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.k_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.k_strm_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.k_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.k_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.k_strm_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.k_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_key_to_mem_U0_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_key_to_mem_U0_U.if_empty_n & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0.ap_idle & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_key_to_mem_U0_U.if_write} start_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_key_to_mem_U0_U.if_empty_n & grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0.ap_idle & ~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_key_to_mem_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_key_to_mem_U0_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.tree_expansion_U0',");
                        end
                    end
                    1: begin //  for dep proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0'
// for dep channel '' info is :
// blk sig is {{ap_done_reg_2 & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0.ap_done & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.ap_done} output_sync}
                        if ((ap_done_reg_2 & grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0.ap_done & ~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.ap_done)) begin
                            $display("//      Blocked by output sync logic with process : 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0'");
                        end
                    end
                    3: begin //  for dep proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0'
// for dep channel '' info is :
// blk sig is {{ap_done_reg_2 & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0.ap_done & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0.ap_done} output_sync}
                        if ((ap_done_reg_2 & grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0.ap_done & ~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0.ap_done)) begin
                            $display("//      Blocked by output sync logic with process : 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0'");
                        end
                    end
                    endcase
                end
                3 : begin // for proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0'
                    case(index2)
                    1: begin //  for dep proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_strm_cp_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0.com_strm_cp_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0.com_strm_cp_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_strm_cp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_strm_cp_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_strm_cp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_strm_cp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_strm_cp_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_strm_cp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel '' info is :
// blk sig is {{ap_done_reg_3 & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0.ap_done & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.ap_done} output_sync}
                        if ((ap_done_reg_3 & grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0.ap_done & ~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0.ap_done)) begin
                            $display("//      Blocked by output sync logic with process : 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0'");
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_com_to_mem_U0_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_com_to_mem_U0_U.if_empty_n & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0.ap_idle & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_com_to_mem_U0_U.if_write} start_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_com_to_mem_U0_U.if_empty_n & grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0.ap_idle & ~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_com_to_mem_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.start_for_com_to_mem_U0_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.seed_gen_U0',");
                        end
                    end
                    2: begin //  for dep proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0'
// for dep channel '' info is :
// blk sig is {{ap_done_reg_3 & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0.ap_done & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0.ap_done} output_sync}
                        if ((ap_done_reg_3 & grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.com_to_mem_U0.ap_done & ~grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0.ap_done)) begin
                            $display("//      Blocked by output sync logic with process : 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ggm_tree_fu_2770.grp_ggm_large_fu_1338.key_to_mem_U0'");
                        end
                    end
                    endcase
                end
                4 : begin // for proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0'
                    case(index2)
                    5: begin //  for dep proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0.grp_expand_seed_Pipeline_PROCESS_CHUNKS_fu_102.r_strm_0_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0.grp_expand_seed_Pipeline_PROCESS_CHUNKS_fu_102.r_strm_0_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_1_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0.grp_expand_seed_Pipeline_PROCESS_CHUNKS_fu_102.r_strm_1_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0.grp_expand_seed_Pipeline_PROCESS_CHUNKS_fu_102.r_strm_1_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_1_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_1_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_build_VOLE_U0_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_build_VOLE_U0_U.if_full_n & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0.ap_start & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_build_VOLE_U0_U.if_read} start_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_build_VOLE_U0_U.if_full_n & grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0.ap_start & ~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_build_VOLE_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_build_VOLE_U0_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0',");
                        end
                    end
                    endcase
                end
                5 : begin // for proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'
                    case(index2)
                    4: begin //  for dep proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.r_strm_0_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.r_strm_0_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_1_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.r_strm_1_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.r_strm_1_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_1_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_1_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.r_strm_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_build_VOLE_U0_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_build_VOLE_U0_U.if_empty_n & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.ap_idle & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_build_VOLE_U0_U.if_write} start_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_build_VOLE_U0_U.if_empty_n & grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.ap_idle & ~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_build_VOLE_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_build_VOLE_U0_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.expand_seed_U0',");
                        end
                    end
                    6: begin //  for dep proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.u_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.u_strm_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.u_strm_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.u_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.u_strm_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.u_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.u_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.u_strm_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.u_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_0_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_0_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_1_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_1_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_1_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_1_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_1_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_2_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_2_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_2_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_2_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_2_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_3_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_3_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_3_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_3_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_3_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_4_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_4_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_4_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_4_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_4_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_5_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_5_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_5_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_5_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_5_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_6_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_6_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_6_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_6_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_6_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_7_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_7_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_7_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_7_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_7_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_8_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_8_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_8_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_8_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_8_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_9_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_9_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_9_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_9_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_9_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_10_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_10_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_10_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_10_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_10_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_11_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_11_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_11_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_11_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_11_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_12_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_12_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_12_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_12_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_12_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_13_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_13_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_13_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_13_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_13_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_14_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_14_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_14_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_14_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_14_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_15_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_15_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_15_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_15_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_15_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_16_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_16_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_16_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_16_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_16_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_17_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_17_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_17_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_17_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_17_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_18_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_18_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_18_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_18_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_18_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_19_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_19_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_19_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_19_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_19_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_20_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_20_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_20_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_20_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_20_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_21_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_21_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_21_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_21_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_21_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_22_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_22_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_22_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_22_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_22_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_23_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_23_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_23_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_23_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_23_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_24_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_24_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_24_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_24_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_24_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_25_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_25_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_25_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_25_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_25_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_26_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_26_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_26_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_26_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_26_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_27_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_27_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_27_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_27_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_27_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_28_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_28_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_28_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_28_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_28_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_29_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_29_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_29_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_29_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_29_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_30_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_30_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_30_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_30_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_30_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_31_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_31_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_31_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_31_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_31_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_32_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_32_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_32_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_32_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_32_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_33_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_33_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_33_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_33_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_33_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_34_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_34_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_34_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_34_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_34_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_35_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_35_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_35_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_35_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_35_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_36_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_36_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_36_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_36_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_36_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_37_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_37_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_37_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_37_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_37_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_38_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_38_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_38_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_38_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_38_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_39_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_39_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_39_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_39_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_39_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_40_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_40_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_40_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_40_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_40_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_41_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_41_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_41_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_41_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_41_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_41_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_41_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_42_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_42_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_42_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_42_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_42_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_43_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_43_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_43_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_43_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_43_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_43_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_43_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_44_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_44_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_44_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_44_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_44_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_45_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_45_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_45_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_45_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_45_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_46_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_46_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_46_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_46_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_46_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_47_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_47_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_47_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_47_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_47_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_48_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_48_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_48_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_48_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_48_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_49_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_49_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_49_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_49_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_49_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_50_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_50_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_50_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_50_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_50_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_51_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_51_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_51_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_51_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_51_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_52_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_52_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_52_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_52_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_52_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_53_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_53_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_53_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_53_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_53_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_54_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_54_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_54_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_54_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_54_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_55_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_55_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_55_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_55_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_55_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_56_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_56_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_56_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_56_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_56_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_57_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_57_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_57_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_57_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_57_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_58_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_58_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_58_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_58_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_58_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_59_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_59_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_59_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_59_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_59_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_60_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_60_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_60_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_60_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_60_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_61_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_61_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_61_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_61_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_61_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_62_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_62_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_62_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_62_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_62_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_63_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_63_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_63_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_63_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_63_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_64_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_64_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_64_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_64_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_64_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_64_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_64_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_64_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_64_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_65_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_65_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_65_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_65_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_65_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_65_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_65_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_65_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_65_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_66_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_66_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_66_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_66_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_66_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_66_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_66_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_66_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_66_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_67_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_67_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_67_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_67_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_67_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_67_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_67_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_67_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_67_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_68_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_68_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_68_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_68_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_68_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_68_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_68_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_68_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_68_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_69_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_69_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_69_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_69_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_69_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_69_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_69_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_69_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_69_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_70_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_70_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_70_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_70_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_70_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_70_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_70_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_70_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_70_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_71_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_71_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_71_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_71_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_71_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_72_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_72_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_72_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_72_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_72_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_73_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_73_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_73_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_73_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_73_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_73_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_73_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_73_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_73_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_74_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_74_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_74_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_74_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_74_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_74_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_74_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_74_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_74_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_75_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_75_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_75_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_75_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_75_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_75_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_75_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_75_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_75_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_76_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_76_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_76_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_76_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_76_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_76_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_76_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_76_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_76_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_77_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_77_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_77_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_77_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_77_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_77_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_77_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_77_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_77_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_78_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_78_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_78_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_78_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_78_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_78_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_78_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_78_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_78_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_79_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_79_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_79_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_79_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_79_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_79_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_79_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_79_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_79_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_80_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_80_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_80_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_80_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_80_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_80_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_80_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_80_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_80_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_81_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_81_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_81_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_81_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_81_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_81_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_81_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_81_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_81_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_82_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_82_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_82_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_82_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_82_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_82_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_82_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_82_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_82_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_83_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_83_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_83_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_83_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_83_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_83_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_83_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_83_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_83_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_84_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_84_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_84_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_84_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_84_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_84_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_84_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_84_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_84_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_85_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_85_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_85_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_85_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_85_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_85_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_85_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_85_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_85_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_86_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_86_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_86_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_86_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_86_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_86_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_86_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_86_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_86_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_87_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_87_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_87_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_87_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_87_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_87_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_87_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_87_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_87_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_88_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_88_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_88_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_88_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_88_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_88_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_88_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_88_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_88_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_89_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_89_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_89_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_89_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_89_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_89_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_89_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_89_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_89_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_90_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_90_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_90_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_90_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_90_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_90_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_90_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_90_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_90_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_91_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_91_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_91_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_91_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_91_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_91_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_91_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_91_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_91_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_92_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_92_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_92_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_92_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_92_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_92_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_92_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_92_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_92_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_93_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_93_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_93_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_93_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_93_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_93_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_93_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_93_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_93_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_94_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_94_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_94_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_94_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_94_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_94_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_94_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_94_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_94_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_95_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_95_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_95_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_95_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_95_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_95_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_95_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_95_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_95_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_96_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_96_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_96_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_96_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_96_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_96_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_96_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_96_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_96_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_97_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_97_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_97_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_97_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_97_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_97_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_97_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_97_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_97_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_98_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_98_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_98_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_98_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_98_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_98_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_98_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_98_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_98_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_99_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_99_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_99_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_99_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_99_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_99_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_99_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_99_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_99_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_100_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_100_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_100_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_100_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_100_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_100_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_100_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_100_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_100_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_101_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_101_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_101_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_101_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_101_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_101_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_101_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_101_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_101_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_102_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_102_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_102_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_102_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_102_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_102_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_102_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_102_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_102_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_103_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_103_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_103_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_103_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_103_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_103_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_103_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_103_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_103_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_104_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_104_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_104_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_104_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_104_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_104_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_104_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_104_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_104_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_105_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_105_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_105_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_105_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_105_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_105_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_105_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_105_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_105_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_106_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_106_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_106_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_106_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_106_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_106_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_106_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_106_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_106_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_107_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_107_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_107_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_107_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_107_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_107_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_107_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_107_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_107_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_108_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_108_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_108_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_108_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_108_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_108_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_108_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_108_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_108_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_109_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_109_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_109_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_109_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_109_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_109_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_109_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_109_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_109_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_110_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_110_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_110_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_110_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_110_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_110_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_110_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_110_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_110_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_111_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_111_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_111_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_111_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_111_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_111_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_111_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_111_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_111_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_112_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_112_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_112_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_112_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_112_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_112_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_112_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_112_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_112_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_113_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_113_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_113_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_113_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_113_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_113_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_113_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_113_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_113_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_114_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_114_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_114_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_114_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_114_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_114_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_114_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_114_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_114_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_115_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_115_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_115_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_115_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_115_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_115_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_115_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_115_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_115_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_116_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_116_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_116_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_116_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_116_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_116_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_116_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_116_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_116_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_117_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_117_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_117_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_117_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_117_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_117_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_117_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_117_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_117_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_118_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_118_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_118_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_118_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_118_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_118_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_118_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_118_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_118_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_119_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_119_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_119_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_119_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_119_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_119_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_119_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_119_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_119_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_120_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_120_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_120_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_120_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_120_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_120_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_120_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_120_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_120_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_121_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_121_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_121_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_121_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_121_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_121_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_121_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_121_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_121_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_122_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_122_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_122_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_122_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_122_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_122_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_122_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_122_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_122_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_123_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_123_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_123_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_123_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_123_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_123_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_123_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_123_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_123_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_124_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_124_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_124_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_124_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_124_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_124_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_124_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_124_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_124_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_125_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_125_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_125_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_125_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_125_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_125_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_125_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_125_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_125_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_126_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_126_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_126_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_126_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_126_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_126_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_126_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_126_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_126_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_127_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_127_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.v_strm_127_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_127_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_127_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_127_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_127_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_127_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_127_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_mem_transfer_U0_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_mem_transfer_U0_U.if_full_n & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.ap_start & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_mem_transfer_U0_U.if_read} start_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_mem_transfer_U0_U.if_full_n & grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.ap_start & ~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_mem_transfer_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_mem_transfer_U0_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0',");
                        end
                    end
                    endcase
                end
                6 : begin // for proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0'
                    case(index2)
                    5: begin //  for dep proc 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.u_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.u_strm_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.u_strm_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.u_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.u_strm_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.u_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.u_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.u_strm_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.u_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_0_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_0_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_1_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_1_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_1_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_1_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_1_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_2_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_2_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_2_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_2_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_2_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_3_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_3_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_3_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_3_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_3_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_4_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_4_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_4_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_4_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_4_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_5_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_5_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_5_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_5_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_5_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_6_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_6_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_6_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_6_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_6_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_7_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_7_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_7_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_7_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_7_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_8_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_8_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_8_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_8_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_8_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_9_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_9_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_9_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_9_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_9_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_10_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_10_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_10_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_10_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_10_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_11_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_11_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_11_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_11_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_11_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_12_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_12_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_12_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_12_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_12_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_13_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_13_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_13_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_13_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_13_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_14_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_14_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_14_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_14_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_14_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_15_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_15_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_15_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_15_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_15_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_16_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_16_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_16_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_16_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_16_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_17_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_17_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_17_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_17_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_17_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_18_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_18_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_18_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_18_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_18_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_19_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_19_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_19_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_19_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_19_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_20_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_20_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_20_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_20_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_20_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_21_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_21_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_21_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_21_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_21_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_22_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_22_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_22_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_22_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_22_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_23_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_23_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_23_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_23_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_23_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_24_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_24_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_24_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_24_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_24_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_25_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_25_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_25_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_25_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_25_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_26_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_26_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_26_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_26_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_26_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_27_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_27_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_27_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_27_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_27_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_28_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_28_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_28_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_28_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_28_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_29_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_29_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_29_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_29_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_29_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_30_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_30_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_30_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_30_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_30_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_31_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_31_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_31_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_31_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_31_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_32_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_32_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_32_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_32_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_32_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_33_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_33_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_33_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_33_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_33_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_34_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_34_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_34_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_34_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_34_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_35_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_35_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_35_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_35_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_35_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_36_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_36_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_36_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_36_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_36_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_37_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_37_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_37_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_37_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_37_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_38_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_38_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_38_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_38_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_38_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_39_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_39_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_39_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_39_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_39_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_40_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_40_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_40_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_40_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_40_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_41_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_41_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_41_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_41_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_41_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_41_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_41_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_42_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_42_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_42_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_42_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_42_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_43_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_43_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_43_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_43_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_43_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_43_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_43_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_44_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_44_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_44_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_44_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_44_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_45_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_45_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_45_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_45_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_45_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_46_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_46_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_46_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_46_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_46_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_47_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_47_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_47_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_47_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_47_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_48_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_48_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_48_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_48_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_48_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_49_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_49_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_49_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_49_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_49_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_50_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_50_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_50_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_50_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_50_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_51_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_51_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_51_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_51_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_51_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_52_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_52_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_52_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_52_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_52_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_53_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_53_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_53_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_53_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_53_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_54_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_54_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_54_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_54_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_54_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_55_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_55_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_55_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_55_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_55_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_56_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_56_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_56_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_56_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_56_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_57_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_57_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_57_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_57_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_57_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_58_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_58_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_58_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_58_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_58_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_59_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_59_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_59_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_59_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_59_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_60_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_60_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_60_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_60_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_60_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_61_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_61_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_61_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_61_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_61_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_62_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_62_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_62_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_62_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_62_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_63_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_63_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_63_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_63_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_63_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_64_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_64_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_64_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_64_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_64_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_64_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_64_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_64_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_64_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_65_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_65_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_65_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_65_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_65_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_65_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_65_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_65_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_65_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_66_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_66_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_66_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_66_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_66_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_66_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_66_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_66_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_66_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_67_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_67_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_67_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_67_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_67_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_67_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_67_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_67_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_67_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_68_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_68_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_68_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_68_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_68_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_68_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_68_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_68_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_68_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_69_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_69_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_69_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_69_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_69_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_69_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_69_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_69_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_69_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_70_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_70_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_70_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_70_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_70_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_70_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_70_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_70_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_70_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_71_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_71_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_71_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_71_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_71_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_72_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_72_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_72_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_72_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_72_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_73_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_73_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_73_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_73_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_73_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_73_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_73_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_73_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_73_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_74_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_74_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_74_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_74_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_74_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_74_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_74_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_74_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_74_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_75_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_75_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_75_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_75_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_75_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_75_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_75_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_75_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_75_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_76_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_76_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_76_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_76_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_76_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_76_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_76_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_76_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_76_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_77_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_77_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_77_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_77_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_77_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_77_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_77_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_77_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_77_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_78_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_78_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_78_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_78_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_78_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_78_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_78_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_78_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_78_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_79_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_79_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_79_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_79_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_79_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_79_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_79_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_79_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_79_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_80_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_80_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_80_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_80_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_80_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_80_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_80_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_80_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_80_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_81_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_81_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_81_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_81_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_81_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_81_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_81_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_81_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_81_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_82_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_82_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_82_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_82_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_82_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_82_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_82_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_82_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_82_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_83_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_83_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_83_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_83_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_83_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_83_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_83_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_83_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_83_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_84_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_84_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_84_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_84_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_84_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_84_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_84_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_84_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_84_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_85_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_85_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_85_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_85_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_85_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_85_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_85_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_85_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_85_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_86_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_86_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_86_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_86_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_86_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_86_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_86_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_86_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_86_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_87_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_87_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_87_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_87_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_87_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_87_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_87_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_87_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_87_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_88_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_88_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_88_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_88_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_88_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_88_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_88_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_88_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_88_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_89_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_89_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_89_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_89_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_89_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_89_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_89_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_89_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_89_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_90_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_90_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_90_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_90_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_90_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_90_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_90_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_90_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_90_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_91_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_91_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_91_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_91_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_91_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_91_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_91_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_91_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_91_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_92_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_92_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_92_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_92_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_92_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_92_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_92_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_92_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_92_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_93_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_93_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_93_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_93_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_93_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_93_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_93_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_93_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_93_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_94_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_94_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_94_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_94_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_94_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_94_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_94_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_94_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_94_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_95_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_95_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_95_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_95_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_95_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_95_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_95_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_95_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_95_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_96_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_96_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_96_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_96_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_96_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_96_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_96_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_96_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_96_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_97_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_97_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_97_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_97_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_97_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_97_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_97_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_97_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_97_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_98_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_98_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_98_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_98_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_98_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_98_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_98_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_98_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_98_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_99_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_99_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_99_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_99_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_99_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_99_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_99_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_99_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_99_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_100_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_100_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_100_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_100_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_100_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_100_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_100_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_100_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_100_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_101_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_101_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_101_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_101_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_101_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_101_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_101_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_101_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_101_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_102_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_102_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_102_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_102_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_102_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_102_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_102_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_102_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_102_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_103_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_103_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_103_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_103_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_103_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_103_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_103_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_103_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_103_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_104_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_104_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_104_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_104_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_104_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_104_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_104_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_104_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_104_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_105_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_105_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_105_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_105_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_105_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_105_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_105_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_105_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_105_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_106_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_106_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_106_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_106_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_106_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_106_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_106_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_106_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_106_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_107_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_107_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_107_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_107_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_107_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_107_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_107_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_107_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_107_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_108_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_108_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_108_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_108_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_108_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_108_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_108_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_108_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_108_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_109_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_109_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_109_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_109_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_109_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_109_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_109_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_109_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_109_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_110_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_110_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_110_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_110_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_110_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_110_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_110_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_110_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_110_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_111_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_111_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_111_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_111_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_111_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_111_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_111_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_111_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_111_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_112_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_112_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_112_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_112_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_112_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_112_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_112_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_112_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_112_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_113_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_113_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_113_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_113_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_113_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_113_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_113_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_113_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_113_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_114_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_114_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_114_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_114_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_114_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_114_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_114_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_114_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_114_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_115_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_115_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_115_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_115_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_115_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_115_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_115_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_115_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_115_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_116_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_116_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_116_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_116_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_116_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_116_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_116_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_116_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_116_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_117_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_117_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_117_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_117_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_117_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_117_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_117_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_117_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_117_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_118_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_118_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_118_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_118_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_118_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_118_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_118_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_118_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_118_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_119_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_119_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_119_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_119_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_119_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_119_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_119_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_119_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_119_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_120_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_120_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_120_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_120_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_120_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_120_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_120_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_120_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_120_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_121_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_121_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_121_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_121_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_121_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_121_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_121_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_121_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_121_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_122_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_122_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_122_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_122_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_122_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_122_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_122_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_122_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_122_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_123_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_123_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_123_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_123_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_123_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_123_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_123_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_123_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_123_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_124_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_124_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_124_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_124_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_124_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_124_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_124_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_124_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_124_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_125_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_125_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_125_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_125_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_125_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_125_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_125_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_125_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_125_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_126_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_126_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_126_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_126_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_126_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_126_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_126_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_126_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_126_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_127_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_127_blk_n data_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.v_strm_127_blk_n)) begin
                            if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_127_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_127_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_127_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_127_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_127_U' read by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.v_strm_127_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_mem_transfer_U0_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_mem_transfer_U0_U.if_empty_n & GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.ap_idle & ~GenerateProof_GenerateProof_inst.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_mem_transfer_U0_U.if_write} start_FIFO}
                        if ((~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_mem_transfer_U0_U.if_empty_n & grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.mem_transfer_U0.ap_idle & ~grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_mem_transfer_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.start_for_mem_transfer_U0_U' written by process 'GenerateProof_GenerateProof.grp_VOLECommit_fu_131.grp_ConvertToVOLE_fu_3305.build_VOLE_U0',");
                        end
                    end
                    endcase
                end
                7 : begin // for proc 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0'
                    case(index2)
                    9: begin //  for dep proc 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.chal2_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.d_strm_cp_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.grp_EvalCircuit_fu_60.grp_EvalCircuit_Pipeline_VITIS_LOOP_100_1_fu_56.d_strm_cp_blk_n data_FIFO} {~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.grp_EvalCircuit_fu_60.grp_EvalCircuit_Pipeline_VITIS_LOOP_107_2_fu_72.d_strm_cp_blk_n data_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.grp_EvalCircuit_fu_60.grp_EvalCircuit_Pipeline_VITIS_LOOP_100_1_fu_56.d_strm_cp_blk_n) | (~grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.grp_EvalCircuit_fu_60.grp_EvalCircuit_Pipeline_VITIS_LOOP_107_2_fu_72.d_strm_cp_blk_n)) begin
                            if (~grp_ProverCircuitEval_fu_148.d_strm_cp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.d_strm_cp_U' written by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.chal2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.d_strm_cp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_ProverCircuitEval_fu_148.d_strm_cp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.d_strm_cp_U' read by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.chal2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.d_strm_cp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.start_for_chal2_U0_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.start_for_chal2_U0_U.if_full_n & GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.ap_start & ~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.real_start & (trans_in_cnt_4 == trans_out_cnt_4) & ~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.start_for_chal2_U0_U.if_read} start_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.start_for_chal2_U0_U.if_full_n & grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.ap_start & ~grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.real_start & (trans_in_cnt_4 == trans_out_cnt_4) & ~grp_ProverCircuitEval_fu_148.start_for_chal2_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.start_for_chal2_U0_U' read by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.chal2_U0',");
                        end
                    end
                    8: begin //  for dep proc 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ToField_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a0_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.grp_EvalCircuit_fu_60.grp_EvalCircuit_Pipeline_VITIS_LOOP_107_2_fu_72.a0_strm_blk_n data_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.grp_EvalCircuit_fu_60.grp_EvalCircuit_Pipeline_VITIS_LOOP_107_2_fu_72.a0_strm_blk_n)) begin
                            if (~grp_ProverCircuitEval_fu_148.a0_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a0_strm_U' written by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ToField_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a0_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_ProverCircuitEval_fu_148.a0_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a0_strm_U' read by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ToField_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a0_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a1_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.grp_EvalCircuit_fu_60.grp_EvalCircuit_Pipeline_VITIS_LOOP_107_2_fu_72.a1_strm_blk_n data_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.grp_EvalCircuit_fu_60.grp_EvalCircuit_Pipeline_VITIS_LOOP_107_2_fu_72.a1_strm_blk_n)) begin
                            if (~grp_ProverCircuitEval_fu_148.a1_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a1_strm_U' written by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ToField_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a1_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_ProverCircuitEval_fu_148.a1_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a1_strm_U' read by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ToField_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a1_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.start_for_ToField_U0_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.start_for_ToField_U0_U.if_full_n & GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.ap_start & ~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.real_start & (trans_in_cnt_4 == trans_out_cnt_4) & ~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.start_for_ToField_U0_U.if_read} start_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.start_for_ToField_U0_U.if_full_n & grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.ap_start & ~grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.real_start & (trans_in_cnt_4 == trans_out_cnt_4) & ~grp_ProverCircuitEval_fu_148.start_for_ToField_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.start_for_ToField_U0_U' read by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ToField_U0',");
                        end
                    end
                    10: begin //  for dep proc 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.aggregate_coef_U0'
// for dep channel '' info is :
// blk sig is {{ap_done_reg_4 & GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.ap_done & ~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.aggregate_coef_U0.ap_done} output_sync}
                        if ((ap_done_reg_4 & grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.ap_done & ~grp_ProverCircuitEval_fu_148.aggregate_coef_U0.ap_done)) begin
                            $display("//      Blocked by output sync logic with process : 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.aggregate_coef_U0'");
                        end
                    end
                    endcase
                end
                8 : begin // for proc 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ToField_U0'
                    case(index2)
                    7: begin //  for dep proc 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a0_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.ToField_U0.a0_strm_blk_n data_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.ToField_U0.a0_strm_blk_n)) begin
                            if (~grp_ProverCircuitEval_fu_148.a0_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a0_strm_U' written by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a0_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_ProverCircuitEval_fu_148.a0_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a0_strm_U' read by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a0_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a1_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.ToField_U0.a1_strm_blk_n data_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.ToField_U0.a1_strm_blk_n)) begin
                            if (~grp_ProverCircuitEval_fu_148.a1_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a1_strm_U' written by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a1_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_ProverCircuitEval_fu_148.a1_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a1_strm_U' read by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a1_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.start_for_ToField_U0_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.start_for_ToField_U0_U.if_empty_n & GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.ToField_U0.ap_idle & ~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.start_for_ToField_U0_U.if_write} start_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.start_for_ToField_U0_U.if_empty_n & grp_ProverCircuitEval_fu_148.ToField_U0.ap_idle & ~grp_ProverCircuitEval_fu_148.start_for_ToField_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.start_for_ToField_U0_U' written by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0',");
                        end
                    end
                    10: begin //  for dep proc 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.aggregate_coef_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.ToField_U0.a_strm_blk_n data_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.ToField_U0.a_strm_blk_n)) begin
                            if (~grp_ProverCircuitEval_fu_148.a_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a_strm_U' written by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.aggregate_coef_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_ProverCircuitEval_fu_148.a_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a_strm_U' read by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.aggregate_coef_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                9 : begin // for proc 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.chal2_U0'
                    case(index2)
                    7: begin //  for dep proc 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.d_strm_cp_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.chal2_U0.d_strm_cp_blk_n data_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.chal2_U0.d_strm_cp_blk_n)) begin
                            if (~grp_ProverCircuitEval_fu_148.d_strm_cp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.d_strm_cp_U' written by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.d_strm_cp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_ProverCircuitEval_fu_148.d_strm_cp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.d_strm_cp_U' read by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.d_strm_cp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.start_for_chal2_U0_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.start_for_chal2_U0_U.if_empty_n & GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.chal2_U0.ap_idle & ~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.start_for_chal2_U0_U.if_write} start_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.start_for_chal2_U0_U.if_empty_n & grp_ProverCircuitEval_fu_148.chal2_U0.ap_idle & ~grp_ProverCircuitEval_fu_148.start_for_chal2_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.start_for_chal2_U0_U' written by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0',");
                        end
                    end
                    10: begin //  for dep proc 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.aggregate_coef_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ch2_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.chal2_U0.grp_shake_extensible_fu_195.ch2_strm_blk_n data_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.chal2_U0.grp_shake_extensible_fu_195.ch2_strm_blk_n)) begin
                            if (~grp_ProverCircuitEval_fu_148.ch2_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ch2_strm_U' written by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.aggregate_coef_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ch2_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_ProverCircuitEval_fu_148.ch2_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ch2_strm_U' read by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.aggregate_coef_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ch2_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                10 : begin // for proc 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.aggregate_coef_U0'
                    case(index2)
                    7: begin //  for dep proc 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.u_mask_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.u_mask_U.if_empty_n & GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.aggregate_coef_U0.ap_idle & ~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.u_mask_U.if_write} TLF_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.u_mask_U.if_empty_n & grp_ProverCircuitEval_fu_148.aggregate_coef_U0.ap_idle & ~grp_ProverCircuitEval_fu_148.u_mask_U.if_write)) begin
                            if (~grp_ProverCircuitEval_fu_148.u_mask_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.u_mask_U' written by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.u_mask_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_ProverCircuitEval_fu_148.u_mask_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.u_mask_U' read by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.u_mask_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.v_mask_U' info is :
// blk sig is {{~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.v_mask_U.if_empty_n & GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.aggregate_coef_U0.ap_idle & ~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.v_mask_U.if_write} TLF_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.v_mask_U.if_empty_n & grp_ProverCircuitEval_fu_148.aggregate_coef_U0.ap_idle & ~grp_ProverCircuitEval_fu_148.v_mask_U.if_write)) begin
                            if (~grp_ProverCircuitEval_fu_148.v_mask_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.v_mask_U' written by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.v_mask_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_ProverCircuitEval_fu_148.v_mask_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.v_mask_U' read by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.v_mask_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel '' info is :
// blk sig is {{ap_done_reg_0 & GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.aggregate_coef_U0.ap_done & ~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.ap_done} output_sync}
                        if ((ap_done_reg_0 & grp_ProverCircuitEval_fu_148.aggregate_coef_U0.ap_done & ~grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0.ap_done)) begin
                            $display("//      Blocked by output sync logic with process : 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ProverCircuitEval_Block_entry_u_0_arg_proc_U0'");
                        end
                    end
                    8: begin //  for dep proc 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ToField_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.aggregate_coef_U0.a_strm_blk_n data_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.aggregate_coef_U0.a_strm_blk_n)) begin
                            if (~grp_ProverCircuitEval_fu_148.a_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a_strm_U' written by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ToField_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_ProverCircuitEval_fu_148.a_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a_strm_U' read by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ToField_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.a_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    9: begin //  for dep proc 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.chal2_U0'
// for dep channel 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ch2_strm_U' info is :
// blk sig is {~GenerateProof_GenerateProof_inst.grp_ProverCircuitEval_fu_148.aggregate_coef_U0.ch2_strm_blk_n data_FIFO}
                        if ((~grp_ProverCircuitEval_fu_148.aggregate_coef_U0.ch2_strm_blk_n)) begin
                            if (~grp_ProverCircuitEval_fu_148.ch2_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ch2_strm_U' written by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.chal2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ch2_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~grp_ProverCircuitEval_fu_148.ch2_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ch2_strm_U' read by process 'GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.chal2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path GenerateProof_GenerateProof.grp_ProverCircuitEval_fu_148.ch2_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
            endcase
        end
    endtask

    // report
    initial begin : report_deadlock
        integer cycle_id;
        integer cycle_comp_id;
        integer record_time;
        wait (dl_reset == 1);
        cycle_id = 1;
        record_time = 0;
        while (1) begin
            @ (negedge dl_clock);
            case (CS_fsm)
                ST_DL_DETECTED: begin
                    cycle_comp_id = 2;
                    if (dl_detect_reg != dl_done_reg && stop_report_path == 1'b0) begin
                        if (dl_done_reg == 'b0) begin
                            print_dl_head;
                            record_time = $time;
                        end
                        print_cycle_start(proc_path(origin), cycle_id);
                        cycle_id = cycle_id + 1;
                    end
                    else begin
                        print_dl_end((cycle_id - 1),record_time);
                        @(negedge dl_clock);
                        @(negedge dl_clock);
                        $finish;
                    end
                end
                ST_DL_REPORT: begin
                    if ((|(dl_in_vec)) & ~(|(dl_in_vec & origin_reg)) & ~(|(reported_proc & dl_in_vec))) begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                        print_cycle_proc_comp(proc_path(dl_in_vec), cycle_comp_id);
                        cycle_comp_id = cycle_comp_id + 1;
                    end
                    else begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                    end
                end
            endcase
        end
    end
 
